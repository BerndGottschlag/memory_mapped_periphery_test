-- Copyright Bernd Gottschlag 2024.
--
-- This source describes Open Hardware and is licensed under the CERN-OHL-W v2
--
-- You may redistribute and modify this documentation and make products using it
-- under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl). This
-- documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED WARRANTY,
-- INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY AND FITNESS FOR A 
-- PARTICULAR PURPOSE. Please see the CERN-OHL-W v2 for applicable conditions.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- This interconnection implements allows a single master node to access two slave nodes

-- Slave 0 (Push buttons) address space: 0x0 to 0x3FF
-- Slave 1 (LEDs) address space: 0x400 to 0x7FF
-- -> i_m0_wb_adr[10] selects the periphery
-- -> a bus error is generated by the intercon if any of i_m0_wb_adr[15 .. 11] is set to 1

entity intercon is
	generic (
		g_WB_DATA_BUS_WIDTH : integer := 8;
		g_M0_WB_ADDRESS_BUS_WIDTH : integer := 16;
		g_S0_WB_ADDRESS_BUS_WIDTH : integer := 10;
		g_S1_WB_ADDRESS_BUS_WIDTH : integer := 10;

		-- address space
		g_S0_ADDRESS_START : integer := 16#0#;
		g_S0_ADDRESS_END : integer := 16#3FF#;

		g_S1_ADDRESS_START : integer := 16#400#;
		g_S1_ADDRESS_END : integer := 16#7FF#
		);
	port (
		-- shared signals
		i_wb_rst : in std_logic;
		i_wb_clk : in std_logic;

		-- master interface (wishbown slave)
		i_m0_wb_dat : in std_logic_vector (g_WB_DATA_BUS_WIDTH - 1 downto 0);
		o_m0_wb_dat : out std_logic_vector (g_WB_DATA_BUS_WIDTH - 1 downto 0);
		i_m0_wb_adr : in std_logic_vector (g_M0_WB_ADDRESS_BUS_WIDTH - 1 downto 0);
		o_m0_wb_ack : out std_logic;
		i_m0_wb_cyc : in std_logic;
		i_m0_wb_stb : in std_logic;
		o_m0_wb_err : out std_logic;
		i_m0_wb_we : in std_logic;

		-- slave 0 interface (wishbown master)
		o_s0_wb_dat : out std_logic_vector (g_WB_DATA_BUS_WIDTH - 1 downto 0);
		i_s0_wb_dat : in std_logic_vector (g_WB_DATA_BUS_WIDTH - 1 downto 0);
		o_s0_wb_adr : out std_logic_vector (g_S0_WB_ADDRESS_BUS_WIDTH - 1 downto 0);
		i_s0_wb_ack : in std_logic;
		o_s0_wb_cyc : out std_logic;
		o_s0_wb_stb : out std_logic;
		i_s0_wb_err : in std_logic;
		o_s0_wb_we : out std_logic;

		-- slave 1 interface (wishbown master)
		o_s1_wb_dat : out std_logic_vector (g_WB_DATA_BUS_WIDTH - 1 downto 0);
		i_s1_wb_dat : in std_logic_vector (g_WB_DATA_BUS_WIDTH - 1 downto 0);
		o_s1_wb_adr : out std_logic_vector (g_S1_WB_ADDRESS_BUS_WIDTH - 1 downto 0);
		i_s1_wb_ack : in std_logic;
		o_s1_wb_cyc : out std_logic;
		o_s1_wb_stb : out std_logic;
		i_s1_wb_err : in std_logic;
		o_s1_wb_we : out std_logic
	);
end;

-- TODO: put inactivation of M0, S0 and S1 in their own functions

architecture rtl of intercon is
	signal r_termination_signaled : std_logic := '0';

	procedure p_DEACTIVATE_M0 (
		signal o_m0_wb_dat : out std_logic_vector (g_WB_DATA_BUS_WIDTH - 1 downto 0);
		signal o_m0_wb_ack : out std_logic;
		signal o_m0_wb_err : out std_logic
	) is
	begin
		o_m0_wb_dat <= std_logic_vector(to_unsigned(0, g_WB_DATA_BUS_WIDTH));
		o_m0_wb_ack <= '0';
		o_m0_wb_err <= '0';
	end p_DEACTIVATE_M0;

	-- Note: there is one deactivation function for each slave as each slave may have a diffrent address width
	procedure p_DEACTIVATE_S0 (
		signal o_s0_wb_dat : out std_logic_vector (g_WB_DATA_BUS_WIDTH - 1 downto 0);
		signal o_s0_wb_adr : out std_logic_vector (g_S0_WB_ADDRESS_BUS_WIDTH - 1 downto 0);
		signal o_s0_wb_cyc : out std_logic;
		signal o_s0_wb_stb : out std_logic;
		signal o_s0_wb_we : out std_logic
	) is
	begin
		o_s0_wb_dat <= std_logic_vector(to_unsigned(0, g_WB_DATA_BUS_WIDTH));
		o_s0_wb_adr <= std_logic_vector(to_unsigned(0, g_S0_WB_ADDRESS_BUS_WIDTH));
		o_s0_wb_cyc <= '0';
		o_s0_wb_stb <= '0';
		o_s0_wb_we <= '0';
	end p_DEACTIVATE_S0;

	procedure p_DEACTIVATE_S1 (
		signal o_s1_wb_dat : out std_logic_vector (g_WB_DATA_BUS_WIDTH - 1 downto 0);
		signal o_s1_wb_adr : out std_logic_vector (g_S1_WB_ADDRESS_BUS_WIDTH - 1 downto 0);
		signal o_s1_wb_cyc : out std_logic;
		signal o_s1_wb_stb : out std_logic;
		signal o_s1_wb_we : out std_logic
	) is
	begin
		o_s1_wb_dat <= std_logic_vector(to_unsigned(0, g_WB_DATA_BUS_WIDTH));
		o_s1_wb_adr <= std_logic_vector(to_unsigned(0, g_S0_WB_ADDRESS_BUS_WIDTH));
		o_s1_wb_cyc <= '0';
		o_s1_wb_stb <= '0';
		o_s1_wb_we <= '0';
	end p_DEACTIVATE_S1;
begin
	p_CONTROL : process (i_wb_clk) is
	begin
		if rising_edge(i_wb_clk) then
			if i_wb_rst = '1' then
					-- set M0 inactive:
					p_DEACTIVATE_M0(o_m0_wb_dat, o_m0_wb_ack, o_m0_wb_err);

					-- set S0 inactive:
					p_DEACTIVATE_S0(o_s0_wb_dat, o_s0_wb_adr, o_s0_wb_cyc, o_s0_wb_stb, o_s0_wb_we);

					-- set S1 inactive:
					p_DEACTIVATE_S1(o_s1_wb_dat, o_s1_wb_adr, o_s1_wb_cyc, o_s1_wb_stb, o_s1_wb_we);

					-- internal signals
					r_termination_signaled <= '0';
			else
				if (i_m0_wb_cyc = '1') AND (i_m0_wb_stb = '1') then
					if (unsigned(i_m0_wb_adr) >= g_S0_ADDRESS_START) AND (unsigned(i_m0_wb_adr) <= g_S0_ADDRESS_END) then
						-- TODO: simplify
						if i_s0_wb_ack = '0' and i_s0_wb_err = '0' and r_termination_signaled = '0' then
							-- connect s0 to m0
							o_s0_wb_dat <= i_m0_wb_dat;
							o_m0_wb_dat <= i_s0_wb_dat;
							o_s0_wb_adr <= i_m0_wb_adr(g_S0_WB_ADDRESS_BUS_WIDTH - 1 downto 0);
							o_s0_wb_cyc <= i_m0_wb_cyc;
							o_s0_wb_stb <= i_m0_wb_stb;
							o_s0_wb_we <= i_m0_wb_we;
						end if;

						if i_s0_wb_ack = '1' or i_s0_wb_err = '1' then
							r_termination_signaled <= '1';

							o_s0_wb_dat <= i_m0_wb_dat;
							o_m0_wb_dat <= i_s0_wb_dat;
							o_m0_wb_ack <= i_s0_wb_ack;
							o_m0_wb_err <= i_s0_wb_err;

							o_s0_wb_cyc <= '0';
							o_s0_wb_stb <= '0';
						end if;
						if r_termination_signaled = '1' then
							-- transaction finished, return to idle state
							p_DEACTIVATE_M0(o_m0_wb_dat, o_m0_wb_ack, o_m0_wb_err);
							p_DEACTIVATE_S0(o_s0_wb_dat, o_s0_wb_adr, o_s0_wb_cyc, o_s0_wb_stb, o_s0_wb_we);
						end if;
					elsif (unsigned(i_m0_wb_adr) >= g_S1_ADDRESS_START) AND (unsigned(i_m0_wb_adr) <= g_S1_ADDRESS_END) then
						-- TODO: simplify
						if i_s1_wb_ack = '0' and i_s1_wb_err = '0' and r_termination_signaled = '0' then
							-- connect s1 to m0
							o_s1_wb_dat <= i_m0_wb_dat;
							o_m0_wb_dat <= i_s1_wb_dat;
							o_s1_wb_adr <= i_m0_wb_adr(g_S0_WB_ADDRESS_BUS_WIDTH - 1 downto 0);
							o_s1_wb_cyc <= i_m0_wb_cyc;
							o_s1_wb_stb <= i_m0_wb_stb;
							o_s1_wb_we <= i_m0_wb_we;
						end if;

						if i_s1_wb_ack = '1' or i_s1_wb_err = '1' then
							r_termination_signaled <= '1';

							o_s1_wb_dat <= i_m0_wb_dat;
							o_m0_wb_dat <= i_s1_wb_dat;
							o_m0_wb_ack <= i_s1_wb_ack;
							o_m0_wb_err <= i_s1_wb_err;

							o_s1_wb_cyc <= '0';
							o_s1_wb_stb <= '0';
						end if;
						if r_termination_signaled = '1' then
							-- transaction finished, return to idle state
							p_DEACTIVATE_M0(o_m0_wb_dat, o_m0_wb_ack, o_m0_wb_err);
							p_DEACTIVATE_S1(o_s1_wb_dat, o_s1_wb_adr, o_s1_wb_cyc, o_s1_wb_stb, o_s1_wb_we);
						end if;
					else
						-- Invalid address, signal the error
						if r_termination_signaled = '0' then
							r_termination_signaled <= '1';
							o_m0_wb_err <= '1';
						else
							o_m0_wb_err <= '0';
						end if;
					end if;
				else
					-- set M0 inactive:
					p_DEACTIVATE_M0(o_m0_wb_dat, o_m0_wb_ack, o_m0_wb_err);

					-- set S0 inactive:
					p_DEACTIVATE_S0(o_s0_wb_dat, o_s0_wb_adr, o_s0_wb_cyc, o_s0_wb_stb, o_s0_wb_we);

					-- set S1 inactive:
					p_DEACTIVATE_S1(o_s1_wb_dat, o_s1_wb_adr, o_s1_wb_cyc, o_s1_wb_stb, o_s1_wb_we);

					-- internal signals
					r_termination_signaled <= '0';
				end if;
			end if;
		end if;
	end process p_CONTROL;
end rtl;
